library verilog;
use verilog.vl_types.all;
entity DigitalFan_vlg_vec_tst is
end DigitalFan_vlg_vec_tst;
